Memristor Random network 
.include ../models/pershin.sub
.model D d
V1 vin gnd sin (0 10.0 1)
Xmem0 vin gnd l0 memristor alpha=0 beta=500000.0 Roff=200000.0 Ron=2000.0 Rinit=200000.0 Vt=0.6
Xmem1 vin n01 l1 memristor alpha=0 beta=500000.0 Roff=200000.0 Ron=2000.0 Rinit=200000.0 Vt=0.6
Xmem2 n01 n11 l2 memristor alpha=0 beta=500000.0 Roff=200000.0 Ron=2000.0 Rinit=200000.0 Vt=0.6
Xmem3 gnd n11 l3 memristor alpha=0 beta=500000.0 Roff=200000.0 Ron=2000.0 Rinit=200000.0 Vt=0.6
.tran 500.0 3 1e-09 uic
.control
run
set wr_vecnames
set wr_singlescale
wrdata /home/ignaciopineyro/MemNet/application/tmp_data/simulation_0_states.csv l0 l1 l2 l3  
wrdata /home/ignaciopineyro/MemNet/application/tmp_data/simulation_0_iv.csv i(v1) vin
quit
.endc
.end
